library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom_y is
    generic (
        DATA_WIDTH : integer := 8;
        ADDR_WIDTH : integer := 4  -- Adjust according to the size of the arrays
    );
    port (
        clk    : in  std_logic;
        addr   : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
        data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
    );
end entity rom_y;

architecture behav of rom_y is
    type rom_type is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);
    signal rom_data : rom_type := (
        "00000001", "00000010", "00000011", "00000100",  -- Example data for X array
        "00000101", "00000110", "00000111", "00001000",
        "00001001", "00001010", "00001011", "00001100",
        "00001101", "00001110", "00001111", "00010000"   -- Example data for Y array
    );
begin
    process(clk)
    begin
        if rising_edge(clk) then
            data <= rom_data(to_integer(unsigned(addr)));
        end if;
    end process;
end architecture behav;

