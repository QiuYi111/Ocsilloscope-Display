library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity rom_y is
    generic (
        DATA_WIDTH : integer := 8;
        ADDR_WIDTH : integer := 14  -- Adjust according to the size of the arrays
    );
    port (
        clk    : in  std_logic;
        addr   : in  std_logic_vector(ADDR_WIDTH-1 downto 0);
        data   : out std_logic_vector(DATA_WIDTH-1 downto 0)
    );
end entity rom_y;

architecture behav of rom_y is
    type rom_type is array (0 to 2**ADDR_WIDTH-1) of std_logic_vector(DATA_WIDTH-1 downto 0);
    signal rom_data : rom_type := (
	 "11101010","11101010","11101000","11101000",
"11100111","11100110","11100101","11100100",
"11100011","11100010","11100001","11100000",
"11011111","11011110","11011101","11011100",
"11011010","11011010","11011000","11011000",
"11010110","11010110","11010100","11010100",
"11010010","11010010","11010000","11001111",
"11001110","11001101","11001100","11001011",
"11001010","11001001","11001000","11000111",
"11000110","11000101","11000100","11000011",
"11000010","11000001","11000000","10111110",
"10111110","10111100","10111100","10111010",
"10111010","10111000","10111000","10110110",
"10110110","10110100","10110100","10110010",
"10110001","10110000","10101111","10101110",
"10101101","10101100","10101011","10101010",
"10101001","10101000","10100111","10100110",
"10100101","10100100","10100010","10100010",
"10100000","10100000","10011110","10011110",
"10011100","10011100","10011010","10011010",
"10011000","10011000","10010110","10010101",
"10010100","10010011","10010010","10010001",
"10010000","10001110","10001101","10001100",
"10001010","10001001","10001000","10000110",
"10000101","10000100","10000010","10000000",
"01111111","01111110","01111100","01111010",
"01111001","01110111","01110101","01110100",
"01110010","01110000","01101110","01101100",
"01101010","01101000","01100110","01100100",
"01100010","01100001","01011111","01011101",
"01011100","01011010","01011000","01010111",
"01010110","01010100","01010010","01010001",
"01010000","01001110","01001101","01001100",
"01001010","01001001","01001000","01000110",
"01000110","01000100","01000011","01000010",
"01000001","01000000","00111111","00111110",
"00111101","00111100","00111011","00111010",
"00111001","00111000","00111000","00110110",
"00110110","00110110","00110100","00110100",
"00110100","00110010","00110010","00110010",
"00110010","00110000","00110000","00110000",
"00110000","00110000","00110000","00110000",
"00110000","00110000","00110000","00110000",
"00110000","00110000","00110000","00110010",
"00110010","00110010","00110011","00110100",
"00110100","00110101","00110110","00110110",
"00111000","00111000","00111001","00111010",
"00111010","00111100","00111100","00111110",
"00111110","01000000","01000000","01000010",
"01000010","01000100","01000100","01000110",
"01000110","01001000","01001001","01001010",
"01001011","01001101","01001111","01010001",
"01010010","01010100","01010101","01010110",
"01010111","01011000","01011010","01011010",
"01011100","01011100","01011110","01011111",
"01100000","01100001","01100010","01100100",
"01100100","01100110","01100110","01101000",
"01101001","01101010","01101011","01101100",
"01101101","01101110","01101111","01110000",
"01110010","01110010","01110100","01110100",
"01110110","01110110","01111000","01111000",
"01111010","01111010","01111100","01111100",
"01111110","01111111","10000000","10000001",
"10000010","10000100","10000101","10000110",
"10001000","10001001","10001011","10001100",
"10001110","10001110","10010000","10010001",
"10010010","10010011","10010100","10010101",
"10010110","10011000","10011001","10011010",
"10011011","10011100","10011101","10011110",
"10011111","10100000","10100010","10100011",
"10100100","10100110","10101000","10101010",
"10101100","10101110","10110000","10110010",
"10110100","10110110","10110110","10110110",
"10110110","10110110","10110100","10110010",
"10110000","10101110","10101101","10101011",
"10101001","10100111","10100101","10100011",
"10100010","10100000","10011111","10011110",
"10011101","10011100","10011011","10011010",
"10011001","10011000","10010111","10010110",
"10010100","10010011","10010010","10010001",
"10010000","10001110","10001101","10001100",
"10001011","10001001","10001000","10000110",
"10000101","10000011","10000010","10000000",
"10000000","01111110","01111101","01111100",
"01111011","01111010","01111010","01111000",
"01111000","01110110","01110110","01110100",
"01110100","01110010","01110010","01110000",
"01110000","01101110","01101110","01101100",
"01101100","01101010","01101010","01101000",
"01101000","01100110","01100101","01100100",
"01100011","01100010","01100000","01100000",
"01011110","01011101","01011100","01011010",
"01011010","01011000","01010111","01010110",
"01010101","01010100","01010010","01010001",
"01010000","01001110","01001101","01001011",
"01001010","01001000","01001000","01000110",
"01000101","01000100","01000011","01000010",
"01000010","01000000","01000000","00111110",
"00111110","00111100","00111100","00111010",
"00111010","00111001","00111000","00111000",
"00110110","00110110","00110110","00110100",
"00110100","00110100","00110011","00110010",
"00110010","00110010","00110010","00110000",
"00110000","00110000","00110000","00110000",
"00110000","00110000","00110000","00110010",
"00110010","00110010","00110010","00110011",
"00110100","00110100","00110100","00110110",
"00110110","00110110","00111000","00111000",
"00111001","00111010","00111010","00111100",
"00111100","00111110","00111110","00111111",
"01000000","01000010","01000010","01000100",
"01000100","01000110","01000111","01001000",
"01001010","01001010","01001100","01001101",
"01001110","01010000","01010001","01010010",
"01010100","01010110","01010111","01011000",
"01011010","01011100","01011101","01011111",
"01100000","01100010","01100100","01100110",
"01101000","01101001","01101011","01101101",
"01101111","01110001","01110010","01110100",
"01110110","01111000","01111001","01111011",
"01111101","01111110","10000000","10000001",
"10000011","10000100","10000110","10000111",
"10001000","10001010","10001011","10001100",
"10001110","10001111","10010000","10010010",
"10010010","10010100","10010101","10010110",
"10010111","10011000","10011010","10011010",
"10011100","10011100","10011110","10011110",
"10100000","10100000","10100010","10100010",
"10100100","10100100","10100110","10100110",
"10101000","10101000","10101010","10101010",
"10101011","10101100","10101101","10101110",
"10101111","10110000","10110001","10110010",
"10110100","10110100","10110110","10110110",
"10110111","10111000","10111001","10111010",
"10111011","10111100","10111101","10111110",
"10111111","11000000","11000001","11000010",
"11000011","11000100","11000101","11000110",
"11000111","11001000","11001001","11001010",
"11001011","11001100","11001101","11001110",
"11001111","11010000","11010001","11010010",
"11010011","11010100","11010101","11010110",
"11010111","11011000","11011001","11011010",
"11011011","11011100","11011101","11011110",
"11011111","11100000","11100001","11100010",
"11100011","11100100","11100101","11100110",
"11100110","11101000","11101000","11101000",
"11101000","11101000","11100111","11100110",
"11100101","11100100","11100010","11100000",
"11011111","11011110","11011100","11011010",
"11011000","11010110","11010100","11010010",
"11010000","11001110","11001100","11001011",
"11001001","11000111","11000101","11000011",
"11000001","11000000","11000000","11000000",
"11000000","11000010","11000100","11000110",
"11001000","11001010","11001100","11001110",
"11010000","11010010","11010100","11010101",
"11010111","11011001","11011011","11011101",
"11011111","11100001","11100010","11100100",
"11100110","11100110","11101000","11101000",
"11101000","11101010","11000111","11000101",
"11000011","11000001","10111111","10111101",
"10111011","10111001","10111000","10110110",
"10110100","10110010","10110000","10101110",
"10101100","10101010","10101000","10101000",
"10100110","10100110","10100100","10100100",
"10100010","10100010","10100000","10100000",
"10011110","10011101","10011100","10011011",
"10011001","10010111","10010101","10010100",
"10010010","10010001","10010000","10001111",
"10001110","10001100","10001100","10001010",
"10001010","10001000","10001000","10000110",
"10000110","10000100","10000100","10000010",
"10000010","10000000","01111111","01111110",
"01111101","01111100","01111011","01111010",
"01111001","01111000","01110111","01110110",
"01110101","01110100","01110011","01110010",
"01110000","01101111","01101110","01101100",
"01101011","01101010","01101000","01100110",
"01100101","01100100","01100010","01100010",
"01100000","01100000","01011110","01011101",
"01011100","01011011","01011010","01011000",
"01011000","01010110","01010110","01010100",
"01010011","01010010","01010001","01010000",
"01001110","01001110","01001100","01001100",
"01001010","01001010","01001000","01001000",
"01000110","01000110","01000110","01000100",
"01000100","01000100","01000100","01000010",
"01000010","01000010","01000010","01000010",
"01000010","01000010","01000010","01000010",
"01000010","01000100","01000100","01000100",
"01000101","01000110","01000110","01000111",
"01001000","01001001","01001010","01001011",
"01001100","01001101","01001110","01001111",
"01010000","01010001","01010010","01010100",
"01010101","01010110","01011000","01011001",
"01011010","01011100","01011101","01011111",
"01100000","01100010","01100100","01100110",
"01100111","01101001","01101011","01101101",
"01101111","01110000","01110010","01110100",
"01110110","01110111","01111001","01111010",
		  others => (others => '0')
		  );
begin
    process(clk)
    begin
        if rising_edge(clk) then
            data <= rom_data(to_integer(unsigned(addr)));
        end if;
    end process;
end architecture behav;

